module Mod3Counter (
    input clk_i,
    input nrst,
    output clk_o
);


    
endmodule
module PC (
    input clk,
    input nrst,
    input [31:0] pc_in,
    output [31:0] pc_out
);


    
endmodule
module LED_test (
    input a,
    input b,
    output c
);
    assign c = a & b;
endmodule
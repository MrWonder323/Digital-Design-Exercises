module Reg_file (
    input clk,
    input addr_in1,
    input addr_in2,
    input addr_in3,
    input data_in3,
    input we3,
    output data_out1,
    output data_out2

);
    
endmodule
module inst_mem (
    input address,
    output [31:0] inst_out
);
    
endmodule